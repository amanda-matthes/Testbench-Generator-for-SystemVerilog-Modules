/*
This is counter with width WIDTH
*/
module counter (
    input wire clk, res_n,
    output reg [WIDTH-1:0] cnt_out
    );                                   
    
    
endmodule

